
package my_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "packet.sv"
    `include "sequence_in.sv"
    `include "monitor.sv"
    `include "driver.sv"
    `include "agent.sv"
    `include "refmod.sv"
    `include "cover_mem.sv"
    `include "scoreboard.sv"
    `include "env.sv"
    `include "tc_sanity.sv"
endpackage

